`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:07:37 01/23/2022 
// Design Name: 
// Module Name:    Dzielnik_1Hz 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Dzielnik_1Hz(
    input in_clock,
    output out_clock
    );
	 
always @(posedge in_clock)
begin 
	
end


endmodule
